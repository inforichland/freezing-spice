library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.common.all;
use work.mem_pkg.all;

entity memory_stage is
    port (mem_d : in  mem_in;
          mem_q : out mem_out);
end entity memory_stage;

architecture Behavioral of memory_stage is
begin  -- architecture Behavioral



end architecture Behavioral;
