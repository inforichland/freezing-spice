library ieee;
use ieee.std_logic_1164.all;

package test_config is

    constant pipeline_tb_test_vector_input_filename : string := "test1.vec";

end package test_config;
